library verilog;
use verilog.vl_types.all;
entity filter_3X3_vlg_tst is
end filter_3X3_vlg_tst;
