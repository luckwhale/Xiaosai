library verilog;
use verilog.vl_types.all;
entity cyclone10lp_routing_wire is
    port(
        datain          : in     vl_logic;
        dataout         : out    vl_logic
    );
end cyclone10lp_routing_wire;
